// CPEN391_Computer.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module CPEN391_Computer (
		output wire [7:0]  hex0_1_export,                   //               hex0_1.export
		output wire [7:0]  hex2_3_export,                   //               hex2_3.export
		output wire [7:0]  hex4_5_export,                   //               hex4_5.export
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //               hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                     .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                     .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                     .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                     .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                     .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                     .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                     .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                     .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                     .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                     .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                     .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                     .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                     .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,     //                     .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,     //                     .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,     //                     .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,     //                     .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,     //                     .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,     //                     .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                     .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                     .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                     .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                     .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                     .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                     .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                     .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                     .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                     .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                     .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                     .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                     .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                     .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                     .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                     .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                     .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                     .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                     .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,    //                     .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,   //                     .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,   //                     .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,    //                     .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                     .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                     .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //                     .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //                     .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //                     .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //                     .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,  //                     .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,  //                     .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,  //                     .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO41,  //                     .hps_io_gpio_inst_GPIO41
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,  //                     .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,  //                     .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,  //                     .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,  //                     .hps_io_gpio_inst_GPIO61
		input  wire        io_acknowledge,                  //                   io.acknowledge
		input  wire        io_irq,                          //                     .irq
		output wire [15:0] io_address,                      //                     .address
		output wire        io_bus_enable,                   //                     .bus_enable
		output wire [1:0]  io_byte_enable,                  //                     .byte_enable
		output wire        io_rw,                           //                     .rw
		output wire [15:0] io_write_data,                   //                     .write_data
		input  wire [15:0] io_read_data,                    //                     .read_data
		output wire [9:0]  leds_export,                     //                 leds.export
		output wire [14:0] memory_mem_a,                    //               memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                     .mem_ba
		output wire        memory_mem_ck,                   //                     .mem_ck
		output wire        memory_mem_ck_n,                 //                     .mem_ck_n
		output wire        memory_mem_cke,                  //                     .mem_cke
		output wire        memory_mem_cs_n,                 //                     .mem_cs_n
		output wire        memory_mem_ras_n,                //                     .mem_ras_n
		output wire        memory_mem_cas_n,                //                     .mem_cas_n
		output wire        memory_mem_we_n,                 //                     .mem_we_n
		output wire        memory_mem_reset_n,              //                     .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                     .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                     .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                     .mem_dqs_n
		output wire        memory_mem_odt,                  //                     .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                     .mem_dm
		input  wire        memory_oct_rzqin,                //                     .oct_rzqin
		input  wire [3:0]  pushbuttons_export,              //          pushbuttons.export
		output wire [12:0] sdram_addr,                      //                sdram.addr
		output wire [1:0]  sdram_ba,                        //                     .ba
		output wire        sdram_cas_n,                     //                     .cas_n
		output wire        sdram_cke,                       //                     .cke
		output wire        sdram_cs_n,                      //                     .cs_n
		inout  wire [15:0] sdram_dq,                        //                     .dq
		output wire [1:0]  sdram_dqm,                       //                     .dqm
		output wire        sdram_ras_n,                     //                     .ras_n
		output wire        sdram_we_n,                      //                     .we_n
		output wire        sdram_clk_clk,                   //            sdram_clk.clk
		input  wire [9:0]  slider_switches_export,          //      slider_switches.export
		input  wire        system_pll_ref_clk_clk,          //   system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset,      // system_pll_ref_reset.reset
		output wire [7:0]  vga_vga_r,                       //                  vga.vga_r
		output wire [7:0]  vga_vga_g,                       //                     .vga_g
		output wire [7:0]  vga_vga_b,                       //                     .vga_b
		output wire        vga_vga_blank_n,                 //                     .vga_blank_n
		output wire        vga_vga_clk,                     //                     .vga_clk
		output wire        vga_vga_hs,                      //                     .vga_hs
		output wire        vga_vga_sync_n,                  //                     .vga_sync_n
		output wire        vga_vga_vs                       //                     .vga_vs
	);

	wire         system_pll_sys_clk_clk;                                             // System_PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, HEX0_1:clk, HEX2_3:clk, HEX4_5:clk, IO_Bridge:clk, Interval_Timer:clk, JTAG_To_FPGA_Bridge:clk_clk, JTAG_To_HPS_Bridge:clk_clk, JTAG_UART_For_ARM0:clk, JTAG_UART_For_ARM1:clk, LEDS:clk, Onchip_SRAM:clk, PushButtons:clk, SDRAM:clk, Slider_Switches:clk, mm_interconnect_0:System_PLL_sys_clk_clk, mm_interconnect_1:System_PLL_sys_clk_clk, renderer_0:clk, rst_controller:clk, rst_controller_003:clk, sysid_qsys_0:clock]
	wire   [1:0] arm_a9_hps_h2f_axi_master_awburst;                                  // ARM_A9_HPS:h2f_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awburst
	wire   [3:0] arm_a9_hps_h2f_axi_master_arlen;                                    // ARM_A9_HPS:h2f_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlen
	wire   [7:0] arm_a9_hps_h2f_axi_master_wstrb;                                    // ARM_A9_HPS:h2f_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wstrb
	wire         arm_a9_hps_h2f_axi_master_wready;                                   // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wready -> ARM_A9_HPS:h2f_WREADY
	wire  [11:0] arm_a9_hps_h2f_axi_master_rid;                                      // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rid -> ARM_A9_HPS:h2f_RID
	wire         arm_a9_hps_h2f_axi_master_rready;                                   // ARM_A9_HPS:h2f_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rready
	wire   [3:0] arm_a9_hps_h2f_axi_master_awlen;                                    // ARM_A9_HPS:h2f_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlen
	wire  [11:0] arm_a9_hps_h2f_axi_master_wid;                                      // ARM_A9_HPS:h2f_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wid
	wire   [3:0] arm_a9_hps_h2f_axi_master_arcache;                                  // ARM_A9_HPS:h2f_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arcache
	wire         arm_a9_hps_h2f_axi_master_wvalid;                                   // ARM_A9_HPS:h2f_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wvalid
	wire  [29:0] arm_a9_hps_h2f_axi_master_araddr;                                   // ARM_A9_HPS:h2f_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_araddr
	wire   [2:0] arm_a9_hps_h2f_axi_master_arprot;                                   // ARM_A9_HPS:h2f_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arprot
	wire   [2:0] arm_a9_hps_h2f_axi_master_awprot;                                   // ARM_A9_HPS:h2f_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awprot
	wire  [63:0] arm_a9_hps_h2f_axi_master_wdata;                                    // ARM_A9_HPS:h2f_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wdata
	wire         arm_a9_hps_h2f_axi_master_arvalid;                                  // ARM_A9_HPS:h2f_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arvalid
	wire   [3:0] arm_a9_hps_h2f_axi_master_awcache;                                  // ARM_A9_HPS:h2f_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awcache
	wire  [11:0] arm_a9_hps_h2f_axi_master_arid;                                     // ARM_A9_HPS:h2f_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arid
	wire   [1:0] arm_a9_hps_h2f_axi_master_arlock;                                   // ARM_A9_HPS:h2f_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlock
	wire   [1:0] arm_a9_hps_h2f_axi_master_awlock;                                   // ARM_A9_HPS:h2f_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlock
	wire  [29:0] arm_a9_hps_h2f_axi_master_awaddr;                                   // ARM_A9_HPS:h2f_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awaddr
	wire   [1:0] arm_a9_hps_h2f_axi_master_bresp;                                    // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bresp -> ARM_A9_HPS:h2f_BRESP
	wire         arm_a9_hps_h2f_axi_master_arready;                                  // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arready -> ARM_A9_HPS:h2f_ARREADY
	wire  [63:0] arm_a9_hps_h2f_axi_master_rdata;                                    // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rdata -> ARM_A9_HPS:h2f_RDATA
	wire         arm_a9_hps_h2f_axi_master_awready;                                  // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awready -> ARM_A9_HPS:h2f_AWREADY
	wire   [1:0] arm_a9_hps_h2f_axi_master_arburst;                                  // ARM_A9_HPS:h2f_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arburst
	wire   [2:0] arm_a9_hps_h2f_axi_master_arsize;                                   // ARM_A9_HPS:h2f_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arsize
	wire         arm_a9_hps_h2f_axi_master_bready;                                   // ARM_A9_HPS:h2f_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bready
	wire         arm_a9_hps_h2f_axi_master_rlast;                                    // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rlast -> ARM_A9_HPS:h2f_RLAST
	wire         arm_a9_hps_h2f_axi_master_wlast;                                    // ARM_A9_HPS:h2f_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wlast
	wire   [1:0] arm_a9_hps_h2f_axi_master_rresp;                                    // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rresp -> ARM_A9_HPS:h2f_RRESP
	wire  [11:0] arm_a9_hps_h2f_axi_master_awid;                                     // ARM_A9_HPS:h2f_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awid
	wire  [11:0] arm_a9_hps_h2f_axi_master_bid;                                      // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bid -> ARM_A9_HPS:h2f_BID
	wire         arm_a9_hps_h2f_axi_master_bvalid;                                   // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bvalid -> ARM_A9_HPS:h2f_BVALID
	wire   [2:0] arm_a9_hps_h2f_axi_master_awsize;                                   // ARM_A9_HPS:h2f_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awsize
	wire         arm_a9_hps_h2f_axi_master_awvalid;                                  // ARM_A9_HPS:h2f_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awvalid
	wire         arm_a9_hps_h2f_axi_master_rvalid;                                   // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rvalid -> ARM_A9_HPS:h2f_RVALID
	wire  [31:0] jtag_to_fpga_bridge_master_readdata;                                // mm_interconnect_0:JTAG_To_FPGA_Bridge_master_readdata -> JTAG_To_FPGA_Bridge:master_readdata
	wire         jtag_to_fpga_bridge_master_waitrequest;                             // mm_interconnect_0:JTAG_To_FPGA_Bridge_master_waitrequest -> JTAG_To_FPGA_Bridge:master_waitrequest
	wire  [31:0] jtag_to_fpga_bridge_master_address;                                 // JTAG_To_FPGA_Bridge:master_address -> mm_interconnect_0:JTAG_To_FPGA_Bridge_master_address
	wire         jtag_to_fpga_bridge_master_read;                                    // JTAG_To_FPGA_Bridge:master_read -> mm_interconnect_0:JTAG_To_FPGA_Bridge_master_read
	wire   [3:0] jtag_to_fpga_bridge_master_byteenable;                              // JTAG_To_FPGA_Bridge:master_byteenable -> mm_interconnect_0:JTAG_To_FPGA_Bridge_master_byteenable
	wire         jtag_to_fpga_bridge_master_readdatavalid;                           // mm_interconnect_0:JTAG_To_FPGA_Bridge_master_readdatavalid -> JTAG_To_FPGA_Bridge:master_readdatavalid
	wire         jtag_to_fpga_bridge_master_write;                                   // JTAG_To_FPGA_Bridge:master_write -> mm_interconnect_0:JTAG_To_FPGA_Bridge_master_write
	wire  [31:0] jtag_to_fpga_bridge_master_writedata;                               // JTAG_To_FPGA_Bridge:master_writedata -> mm_interconnect_0:JTAG_To_FPGA_Bridge_master_writedata
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;                               // ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awburst
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;                                 // ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlen
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;                                 // ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	wire         arm_a9_hps_h2f_lw_axi_master_wready;                                // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_rid;                                   // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	wire         arm_a9_hps_h2f_lw_axi_master_rready;                                // ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rready
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;                                 // ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlen
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_wid;                                   // ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;                               // ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arcache
	wire         arm_a9_hps_h2f_lw_axi_master_wvalid;                                // ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;                                // ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_araddr
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;                                // ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arprot
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;                                // ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awprot
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;                                 // ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wdata
	wire         arm_a9_hps_h2f_lw_axi_master_arvalid;                               // ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	wire   [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;                               // ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awcache
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_arid;                                  // ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arid
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;                                // ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlock
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;                                // ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlock
	wire  [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;                                // ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;                                 // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	wire         arm_a9_hps_h2f_lw_axi_master_arready;                               // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	wire  [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;                                 // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	wire         arm_a9_hps_h2f_lw_axi_master_awready;                               // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;                               // ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arburst
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;                                // ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arsize
	wire         arm_a9_hps_h2f_lw_axi_master_bready;                                // ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bready
	wire         arm_a9_hps_h2f_lw_axi_master_rlast;                                 // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	wire         arm_a9_hps_h2f_lw_axi_master_wlast;                                 // ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wlast
	wire   [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;                                 // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_awid;                                  // ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awid
	wire  [11:0] arm_a9_hps_h2f_lw_axi_master_bid;                                   // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	wire         arm_a9_hps_h2f_lw_axi_master_bvalid;                                // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	wire   [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;                                // ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awsize
	wire         arm_a9_hps_h2f_lw_axi_master_awvalid;                               // ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	wire         arm_a9_hps_h2f_lw_axi_master_rvalid;                                // mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	wire         mm_interconnect_0_sdram_s1_chipselect;                              // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                             // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                 // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                    // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                              // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                           // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                   // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                               // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_onchip_sram_s1_chipselect;                        // mm_interconnect_0:Onchip_SRAM_s1_chipselect -> Onchip_SRAM:chipselect
	wire  [31:0] mm_interconnect_0_onchip_sram_s1_readdata;                          // Onchip_SRAM:readdata -> mm_interconnect_0:Onchip_SRAM_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_sram_s1_address;                           // mm_interconnect_0:Onchip_SRAM_s1_address -> Onchip_SRAM:address
	wire   [3:0] mm_interconnect_0_onchip_sram_s1_byteenable;                        // mm_interconnect_0:Onchip_SRAM_s1_byteenable -> Onchip_SRAM:byteenable
	wire         mm_interconnect_0_onchip_sram_s1_write;                             // mm_interconnect_0:Onchip_SRAM_s1_write -> Onchip_SRAM:write
	wire  [31:0] mm_interconnect_0_onchip_sram_s1_writedata;                         // mm_interconnect_0:Onchip_SRAM_s1_writedata -> Onchip_SRAM:writedata
	wire         mm_interconnect_0_onchip_sram_s1_clken;                             // mm_interconnect_0:Onchip_SRAM_s1_clken -> Onchip_SRAM:clken
	wire         mm_interconnect_0_io_bridge_avalon_slave_chipselect;                // mm_interconnect_0:IO_Bridge_avalon_slave_chipselect -> IO_Bridge:avalon_chipselect
	wire  [15:0] mm_interconnect_0_io_bridge_avalon_slave_readdata;                  // IO_Bridge:avalon_readdata -> mm_interconnect_0:IO_Bridge_avalon_slave_readdata
	wire         mm_interconnect_0_io_bridge_avalon_slave_waitrequest;               // IO_Bridge:avalon_waitrequest -> mm_interconnect_0:IO_Bridge_avalon_slave_waitrequest
	wire  [14:0] mm_interconnect_0_io_bridge_avalon_slave_address;                   // mm_interconnect_0:IO_Bridge_avalon_slave_address -> IO_Bridge:avalon_address
	wire         mm_interconnect_0_io_bridge_avalon_slave_read;                      // mm_interconnect_0:IO_Bridge_avalon_slave_read -> IO_Bridge:avalon_read
	wire   [1:0] mm_interconnect_0_io_bridge_avalon_slave_byteenable;                // mm_interconnect_0:IO_Bridge_avalon_slave_byteenable -> IO_Bridge:avalon_byteenable
	wire         mm_interconnect_0_io_bridge_avalon_slave_write;                     // mm_interconnect_0:IO_Bridge_avalon_slave_write -> IO_Bridge:avalon_write
	wire  [15:0] mm_interconnect_0_io_bridge_avalon_slave_writedata;                 // mm_interconnect_0:IO_Bridge_avalon_slave_writedata -> IO_Bridge:avalon_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;              // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;               // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire         mm_interconnect_0_leds_s1_chipselect;                               // mm_interconnect_0:LEDS_s1_chipselect -> LEDS:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                 // LEDS:readdata -> mm_interconnect_0:LEDS_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                  // mm_interconnect_0:LEDS_s1_address -> LEDS:address
	wire         mm_interconnect_0_leds_s1_write;                                    // mm_interconnect_0:LEDS_s1_write -> LEDS:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                // mm_interconnect_0:LEDS_s1_writedata -> LEDS:writedata
	wire         mm_interconnect_0_hex4_5_s1_chipselect;                             // mm_interconnect_0:HEX4_5_s1_chipselect -> HEX4_5:chipselect
	wire  [31:0] mm_interconnect_0_hex4_5_s1_readdata;                               // HEX4_5:readdata -> mm_interconnect_0:HEX4_5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex4_5_s1_address;                                // mm_interconnect_0:HEX4_5_s1_address -> HEX4_5:address
	wire         mm_interconnect_0_hex4_5_s1_write;                                  // mm_interconnect_0:HEX4_5_s1_write -> HEX4_5:write_n
	wire  [31:0] mm_interconnect_0_hex4_5_s1_writedata;                              // mm_interconnect_0:HEX4_5_s1_writedata -> HEX4_5:writedata
	wire         mm_interconnect_0_hex2_3_s1_chipselect;                             // mm_interconnect_0:HEX2_3_s1_chipselect -> HEX2_3:chipselect
	wire  [31:0] mm_interconnect_0_hex2_3_s1_readdata;                               // HEX2_3:readdata -> mm_interconnect_0:HEX2_3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex2_3_s1_address;                                // mm_interconnect_0:HEX2_3_s1_address -> HEX2_3:address
	wire         mm_interconnect_0_hex2_3_s1_write;                                  // mm_interconnect_0:HEX2_3_s1_write -> HEX2_3:write_n
	wire  [31:0] mm_interconnect_0_hex2_3_s1_writedata;                              // mm_interconnect_0:HEX2_3_s1_writedata -> HEX2_3:writedata
	wire         mm_interconnect_0_hex0_1_s1_chipselect;                             // mm_interconnect_0:HEX0_1_s1_chipselect -> HEX0_1:chipselect
	wire  [31:0] mm_interconnect_0_hex0_1_s1_readdata;                               // HEX0_1:readdata -> mm_interconnect_0:HEX0_1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_1_s1_address;                                // mm_interconnect_0:HEX0_1_s1_address -> HEX0_1:address
	wire         mm_interconnect_0_hex0_1_s1_write;                                  // mm_interconnect_0:HEX0_1_s1_write -> HEX0_1:write_n
	wire  [31:0] mm_interconnect_0_hex0_1_s1_writedata;                              // mm_interconnect_0:HEX0_1_s1_writedata -> HEX0_1:writedata
	wire  [31:0] mm_interconnect_0_slider_switches_s1_readdata;                      // Slider_Switches:readdata -> mm_interconnect_0:Slider_Switches_s1_readdata
	wire   [1:0] mm_interconnect_0_slider_switches_s1_address;                       // mm_interconnect_0:Slider_Switches_s1_address -> Slider_Switches:address
	wire         mm_interconnect_0_pushbuttons_s1_chipselect;                        // mm_interconnect_0:PushButtons_s1_chipselect -> PushButtons:chipselect
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_readdata;                          // PushButtons:readdata -> mm_interconnect_0:PushButtons_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbuttons_s1_address;                           // mm_interconnect_0:PushButtons_s1_address -> PushButtons:address
	wire         mm_interconnect_0_pushbuttons_s1_write;                             // mm_interconnect_0:PushButtons_s1_write -> PushButtons:write_n
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_writedata;                         // mm_interconnect_0:PushButtons_s1_writedata -> PushButtons:writedata
	wire         mm_interconnect_0_interval_timer_s1_chipselect;                     // mm_interconnect_0:Interval_Timer_s1_chipselect -> Interval_Timer:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_s1_readdata;                       // Interval_Timer:readdata -> mm_interconnect_0:Interval_Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_s1_address;                        // mm_interconnect_0:Interval_Timer_s1_address -> Interval_Timer:address
	wire         mm_interconnect_0_interval_timer_s1_write;                          // mm_interconnect_0:Interval_Timer_s1_write -> Interval_Timer:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_s1_writedata;                      // mm_interconnect_0:Interval_Timer_s1_writedata -> Interval_Timer:writedata
	wire  [31:0] mm_interconnect_0_renderer_0_slave_readdata;                        // renderer_0:slave_readdata -> mm_interconnect_0:renderer_0_slave_readdata
	wire         mm_interconnect_0_renderer_0_slave_waitrequest;                     // renderer_0:slave_waitrequest -> mm_interconnect_0:renderer_0_slave_waitrequest
	wire   [3:0] mm_interconnect_0_renderer_0_slave_address;                         // mm_interconnect_0:renderer_0_slave_address -> renderer_0:slave_address
	wire         mm_interconnect_0_renderer_0_slave_read;                            // mm_interconnect_0:renderer_0_slave_read -> renderer_0:slave_read
	wire         mm_interconnect_0_renderer_0_slave_write;                           // mm_interconnect_0:renderer_0_slave_write -> renderer_0:slave_write
	wire  [31:0] mm_interconnect_0_renderer_0_slave_writedata;                       // mm_interconnect_0:renderer_0_slave_writedata -> renderer_0:slave_writedata
	wire         mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_UART_For_ARM0_avalon_jtag_slave_chipselect -> JTAG_UART_For_ARM0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_readdata;    // JTAG_UART_For_ARM0:av_readdata -> mm_interconnect_0:JTAG_UART_For_ARM0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_waitrequest; // JTAG_UART_For_ARM0:av_waitrequest -> mm_interconnect_0:JTAG_UART_For_ARM0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_UART_For_ARM0_avalon_jtag_slave_address -> JTAG_UART_For_ARM0:av_address
	wire         mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_UART_For_ARM0_avalon_jtag_slave_read -> JTAG_UART_For_ARM0:av_read_n
	wire         mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_UART_For_ARM0_avalon_jtag_slave_write -> JTAG_UART_For_ARM0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_UART_For_ARM0_avalon_jtag_slave_writedata -> JTAG_UART_For_ARM0:av_writedata
	wire         mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_UART_For_ARM1_avalon_jtag_slave_chipselect -> JTAG_UART_For_ARM1:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_readdata;    // JTAG_UART_For_ARM1:av_readdata -> mm_interconnect_0:JTAG_UART_For_ARM1_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_waitrequest; // JTAG_UART_For_ARM1:av_waitrequest -> mm_interconnect_0:JTAG_UART_For_ARM1_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_UART_For_ARM1_avalon_jtag_slave_address -> JTAG_UART_For_ARM1:av_address
	wire         mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_UART_For_ARM1_avalon_jtag_slave_read -> JTAG_UART_For_ARM1:av_read_n
	wire         mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_UART_For_ARM1_avalon_jtag_slave_write -> JTAG_UART_For_ARM1:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_UART_For_ARM1_avalon_jtag_slave_writedata -> JTAG_UART_For_ARM1:av_writedata
	wire  [31:0] jtag_to_hps_bridge_master_readdata;                                 // mm_interconnect_1:JTAG_To_HPS_Bridge_master_readdata -> JTAG_To_HPS_Bridge:master_readdata
	wire         jtag_to_hps_bridge_master_waitrequest;                              // mm_interconnect_1:JTAG_To_HPS_Bridge_master_waitrequest -> JTAG_To_HPS_Bridge:master_waitrequest
	wire  [31:0] jtag_to_hps_bridge_master_address;                                  // JTAG_To_HPS_Bridge:master_address -> mm_interconnect_1:JTAG_To_HPS_Bridge_master_address
	wire         jtag_to_hps_bridge_master_read;                                     // JTAG_To_HPS_Bridge:master_read -> mm_interconnect_1:JTAG_To_HPS_Bridge_master_read
	wire   [3:0] jtag_to_hps_bridge_master_byteenable;                               // JTAG_To_HPS_Bridge:master_byteenable -> mm_interconnect_1:JTAG_To_HPS_Bridge_master_byteenable
	wire         jtag_to_hps_bridge_master_readdatavalid;                            // mm_interconnect_1:JTAG_To_HPS_Bridge_master_readdatavalid -> JTAG_To_HPS_Bridge:master_readdatavalid
	wire         jtag_to_hps_bridge_master_write;                                    // JTAG_To_HPS_Bridge:master_write -> mm_interconnect_1:JTAG_To_HPS_Bridge_master_write
	wire  [31:0] jtag_to_hps_bridge_master_writedata;                                // JTAG_To_HPS_Bridge:master_writedata -> mm_interconnect_1:JTAG_To_HPS_Bridge_master_writedata
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst;                 // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awburst -> ARM_A9_HPS:f2h_AWBURST
	wire   [4:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awuser -> ARM_A9_HPS:f2h_AWUSER
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen;                   // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arlen -> ARM_A9_HPS:f2h_ARLEN
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb;                   // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wstrb -> ARM_A9_HPS:f2h_WSTRB
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready;                  // ARM_A9_HPS:f2h_WREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wready
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid;                     // ARM_A9_HPS:f2h_RID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rid
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rready -> ARM_A9_HPS:f2h_RREADY
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen;                   // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awlen -> ARM_A9_HPS:f2h_AWLEN
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid;                     // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wid -> ARM_A9_HPS:f2h_WID
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache;                 // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arcache -> ARM_A9_HPS:f2h_ARCACHE
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wvalid -> ARM_A9_HPS:f2h_WVALID
	wire  [31:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_araddr -> ARM_A9_HPS:f2h_ARADDR
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arprot -> ARM_A9_HPS:f2h_ARPROT
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awprot -> ARM_A9_HPS:f2h_AWPROT
	wire  [63:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata;                   // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wdata -> ARM_A9_HPS:f2h_WDATA
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid;                 // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arvalid -> ARM_A9_HPS:f2h_ARVALID
	wire   [3:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache;                 // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awcache -> ARM_A9_HPS:f2h_AWCACHE
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid;                    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arid -> ARM_A9_HPS:f2h_ARID
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arlock -> ARM_A9_HPS:f2h_ARLOCK
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awlock -> ARM_A9_HPS:f2h_AWLOCK
	wire  [31:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awaddr -> ARM_A9_HPS:f2h_AWADDR
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp;                   // ARM_A9_HPS:f2h_BRESP -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bresp
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready;                 // ARM_A9_HPS:f2h_ARREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arready
	wire  [63:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata;                   // ARM_A9_HPS:f2h_RDATA -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rdata
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready;                 // ARM_A9_HPS:f2h_AWREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awready
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst;                 // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arburst -> ARM_A9_HPS:f2h_ARBURST
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arsize -> ARM_A9_HPS:f2h_ARSIZE
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bready -> ARM_A9_HPS:f2h_BREADY
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast;                   // ARM_A9_HPS:f2h_RLAST -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rlast
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast;                   // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wlast -> ARM_A9_HPS:f2h_WLAST
	wire   [1:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp;                   // ARM_A9_HPS:f2h_RRESP -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rresp
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid;                    // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awid -> ARM_A9_HPS:f2h_AWID
	wire   [7:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid;                     // ARM_A9_HPS:f2h_BID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bid
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid;                  // ARM_A9_HPS:f2h_BVALID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bvalid
	wire   [2:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awsize -> ARM_A9_HPS:f2h_AWSIZE
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid;                 // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awvalid -> ARM_A9_HPS:f2h_AWVALID
	wire   [4:0] mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser;                  // mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_aruser -> ARM_A9_HPS:f2h_ARUSER
	wire         mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid;                  // ARM_A9_HPS:f2h_RVALID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rvalid
	wire         irq_mapper_receiver0_irq;                                           // IO_Bridge:avalon_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                           // PushButtons:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                           // JTAG_UART_For_ARM0:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                           // Interval_Timer:irq -> irq_mapper:receiver3_irq
	wire  [31:0] arm_a9_hps_f2h_irq0_irq;                                            // irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	wire         irq_mapper_001_receiver0_irq;                                       // JTAG_UART_For_ARM1:av_irq -> irq_mapper_001:receiver0_irq
	wire  [31:0] arm_a9_hps_f2h_irq1_irq;                                            // irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [HEX0_1:reset_n, HEX2_3:reset_n, HEX4_5:reset_n, IO_Bridge:reset, Interval_Timer:reset_n, JTAG_UART_For_ARM0:rst_n, JTAG_UART_For_ARM1:rst_n, LEDS:reset_n, Onchip_SRAM:reset, PushButtons:reset_n, SDRAM:reset_n, Slider_Switches:reset_n, mm_interconnect_0:JTAG_To_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:SDRAM_reset_reset_bridge_in_reset_reset, mm_interconnect_1:JTAG_To_HPS_Bridge_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:JTAG_To_HPS_Bridge_master_translator_reset_reset_bridge_in_reset_reset, renderer_0:rst_n, rst_translator:in_reset, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                 // rst_controller:reset_req -> [Onchip_SRAM:reset_req, rst_translator:reset_req_in]
	wire         arm_a9_hps_h2f_reset_reset;                                         // ARM_A9_HPS:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	wire         system_pll_reset_source_reset;                                      // System_PLL:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> JTAG_To_FPGA_Bridge:clk_reset_reset
	wire         rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> JTAG_To_HPS_Bridge:clk_reset_reset
	wire         rst_controller_003_reset_out_reset;                                 // rst_controller_003:reset_out -> [mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]

	CPEN391_Computer_ARM_A9_HPS #(
		.F2S_Width (2),
		.S2F_Width (2)
	) arm_a9_hps (
		.h2f_mpu_eventi           (),                                                   //    h2f_mpu_events.eventi
		.h2f_mpu_evento           (),                                                   //                  .evento
		.h2f_mpu_standbywfe       (),                                                   //                  .standbywfe
		.h2f_mpu_standbywfi       (),                                                   //                  .standbywfi
		.mem_a                    (memory_mem_a),                                       //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                      //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                      //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                    //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                     //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                    //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                   //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                   //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                    //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                 //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                      //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                     //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                   //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                     //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                      //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                   //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),                    //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                      //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                      //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                      //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                      //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                      //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                      //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                       //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),                    //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),                    //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),                    //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                      //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                      //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                      //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),                        //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),                        //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),                        //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),                        //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),                        //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),                        //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                        //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                         //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                         //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                        //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                         //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                         //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                         //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                         //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                         //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                         //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                         //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                         //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                         //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                         //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                        //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                        //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                        //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                        //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),                       //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),                      //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),                      //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),                       //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                        //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                        //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                        //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                        //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),                        //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),                        //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),                     //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),                     //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),                     //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_io_hps_io_gpio_inst_GPIO41),                     //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),                     //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),                     //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),                     //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),                     //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (arm_a9_hps_h2f_reset_reset),                         //         h2f_reset.reset_n
		.h2f_axi_clk              (system_pll_sys_clk_clk),                             //     h2f_axi_clock.clk
		.h2f_AWID                 (arm_a9_hps_h2f_axi_master_awid),                     //    h2f_axi_master.awid
		.h2f_AWADDR               (arm_a9_hps_h2f_axi_master_awaddr),                   //                  .awaddr
		.h2f_AWLEN                (arm_a9_hps_h2f_axi_master_awlen),                    //                  .awlen
		.h2f_AWSIZE               (arm_a9_hps_h2f_axi_master_awsize),                   //                  .awsize
		.h2f_AWBURST              (arm_a9_hps_h2f_axi_master_awburst),                  //                  .awburst
		.h2f_AWLOCK               (arm_a9_hps_h2f_axi_master_awlock),                   //                  .awlock
		.h2f_AWCACHE              (arm_a9_hps_h2f_axi_master_awcache),                  //                  .awcache
		.h2f_AWPROT               (arm_a9_hps_h2f_axi_master_awprot),                   //                  .awprot
		.h2f_AWVALID              (arm_a9_hps_h2f_axi_master_awvalid),                  //                  .awvalid
		.h2f_AWREADY              (arm_a9_hps_h2f_axi_master_awready),                  //                  .awready
		.h2f_WID                  (arm_a9_hps_h2f_axi_master_wid),                      //                  .wid
		.h2f_WDATA                (arm_a9_hps_h2f_axi_master_wdata),                    //                  .wdata
		.h2f_WSTRB                (arm_a9_hps_h2f_axi_master_wstrb),                    //                  .wstrb
		.h2f_WLAST                (arm_a9_hps_h2f_axi_master_wlast),                    //                  .wlast
		.h2f_WVALID               (arm_a9_hps_h2f_axi_master_wvalid),                   //                  .wvalid
		.h2f_WREADY               (arm_a9_hps_h2f_axi_master_wready),                   //                  .wready
		.h2f_BID                  (arm_a9_hps_h2f_axi_master_bid),                      //                  .bid
		.h2f_BRESP                (arm_a9_hps_h2f_axi_master_bresp),                    //                  .bresp
		.h2f_BVALID               (arm_a9_hps_h2f_axi_master_bvalid),                   //                  .bvalid
		.h2f_BREADY               (arm_a9_hps_h2f_axi_master_bready),                   //                  .bready
		.h2f_ARID                 (arm_a9_hps_h2f_axi_master_arid),                     //                  .arid
		.h2f_ARADDR               (arm_a9_hps_h2f_axi_master_araddr),                   //                  .araddr
		.h2f_ARLEN                (arm_a9_hps_h2f_axi_master_arlen),                    //                  .arlen
		.h2f_ARSIZE               (arm_a9_hps_h2f_axi_master_arsize),                   //                  .arsize
		.h2f_ARBURST              (arm_a9_hps_h2f_axi_master_arburst),                  //                  .arburst
		.h2f_ARLOCK               (arm_a9_hps_h2f_axi_master_arlock),                   //                  .arlock
		.h2f_ARCACHE              (arm_a9_hps_h2f_axi_master_arcache),                  //                  .arcache
		.h2f_ARPROT               (arm_a9_hps_h2f_axi_master_arprot),                   //                  .arprot
		.h2f_ARVALID              (arm_a9_hps_h2f_axi_master_arvalid),                  //                  .arvalid
		.h2f_ARREADY              (arm_a9_hps_h2f_axi_master_arready),                  //                  .arready
		.h2f_RID                  (arm_a9_hps_h2f_axi_master_rid),                      //                  .rid
		.h2f_RDATA                (arm_a9_hps_h2f_axi_master_rdata),                    //                  .rdata
		.h2f_RRESP                (arm_a9_hps_h2f_axi_master_rresp),                    //                  .rresp
		.h2f_RLAST                (arm_a9_hps_h2f_axi_master_rlast),                    //                  .rlast
		.h2f_RVALID               (arm_a9_hps_h2f_axi_master_rvalid),                   //                  .rvalid
		.h2f_RREADY               (arm_a9_hps_h2f_axi_master_rready),                   //                  .rready
		.f2h_axi_clk              (system_pll_sys_clk_clk),                             //     f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr),  //                  .awaddr
		.f2h_AWLEN                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen),   //                  .awlen
		.f2h_AWSIZE               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize),  //                  .awsize
		.f2h_AWBURST              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst), //                  .awburst
		.f2h_AWLOCK               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock),  //                  .awlock
		.f2h_AWCACHE              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache), //                  .awcache
		.f2h_AWPROT               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot),  //                  .awprot
		.f2h_AWVALID              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid), //                  .awvalid
		.f2h_AWREADY              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready), //                  .awready
		.f2h_AWUSER               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser),  //                  .awuser
		.f2h_WID                  (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid),     //                  .wid
		.f2h_WDATA                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata),   //                  .wdata
		.f2h_WSTRB                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb),   //                  .wstrb
		.f2h_WLAST                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast),   //                  .wlast
		.f2h_WVALID               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid),  //                  .wvalid
		.f2h_WREADY               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready),  //                  .wready
		.f2h_BID                  (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid),     //                  .bid
		.f2h_BRESP                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp),   //                  .bresp
		.f2h_BVALID               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid),  //                  .bvalid
		.f2h_BREADY               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready),  //                  .bready
		.f2h_ARID                 (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid),    //                  .arid
		.f2h_ARADDR               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr),  //                  .araddr
		.f2h_ARLEN                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen),   //                  .arlen
		.f2h_ARSIZE               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize),  //                  .arsize
		.f2h_ARBURST              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst), //                  .arburst
		.f2h_ARLOCK               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock),  //                  .arlock
		.f2h_ARCACHE              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache), //                  .arcache
		.f2h_ARPROT               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot),  //                  .arprot
		.f2h_ARVALID              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid), //                  .arvalid
		.f2h_ARREADY              (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready), //                  .arready
		.f2h_ARUSER               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser),  //                  .aruser
		.f2h_RID                  (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid),     //                  .rid
		.f2h_RDATA                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata),   //                  .rdata
		.f2h_RRESP                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp),   //                  .rresp
		.f2h_RLAST                (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast),   //                  .rlast
		.f2h_RVALID               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid),  //                  .rvalid
		.f2h_RREADY               (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready),  //                  .rready
		.h2f_lw_axi_clk           (system_pll_sys_clk_clk),                             //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (arm_a9_hps_h2f_lw_axi_master_awid),                  // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (arm_a9_hps_h2f_lw_axi_master_awaddr),                //                  .awaddr
		.h2f_lw_AWLEN             (arm_a9_hps_h2f_lw_axi_master_awlen),                 //                  .awlen
		.h2f_lw_AWSIZE            (arm_a9_hps_h2f_lw_axi_master_awsize),                //                  .awsize
		.h2f_lw_AWBURST           (arm_a9_hps_h2f_lw_axi_master_awburst),               //                  .awburst
		.h2f_lw_AWLOCK            (arm_a9_hps_h2f_lw_axi_master_awlock),                //                  .awlock
		.h2f_lw_AWCACHE           (arm_a9_hps_h2f_lw_axi_master_awcache),               //                  .awcache
		.h2f_lw_AWPROT            (arm_a9_hps_h2f_lw_axi_master_awprot),                //                  .awprot
		.h2f_lw_AWVALID           (arm_a9_hps_h2f_lw_axi_master_awvalid),               //                  .awvalid
		.h2f_lw_AWREADY           (arm_a9_hps_h2f_lw_axi_master_awready),               //                  .awready
		.h2f_lw_WID               (arm_a9_hps_h2f_lw_axi_master_wid),                   //                  .wid
		.h2f_lw_WDATA             (arm_a9_hps_h2f_lw_axi_master_wdata),                 //                  .wdata
		.h2f_lw_WSTRB             (arm_a9_hps_h2f_lw_axi_master_wstrb),                 //                  .wstrb
		.h2f_lw_WLAST             (arm_a9_hps_h2f_lw_axi_master_wlast),                 //                  .wlast
		.h2f_lw_WVALID            (arm_a9_hps_h2f_lw_axi_master_wvalid),                //                  .wvalid
		.h2f_lw_WREADY            (arm_a9_hps_h2f_lw_axi_master_wready),                //                  .wready
		.h2f_lw_BID               (arm_a9_hps_h2f_lw_axi_master_bid),                   //                  .bid
		.h2f_lw_BRESP             (arm_a9_hps_h2f_lw_axi_master_bresp),                 //                  .bresp
		.h2f_lw_BVALID            (arm_a9_hps_h2f_lw_axi_master_bvalid),                //                  .bvalid
		.h2f_lw_BREADY            (arm_a9_hps_h2f_lw_axi_master_bready),                //                  .bready
		.h2f_lw_ARID              (arm_a9_hps_h2f_lw_axi_master_arid),                  //                  .arid
		.h2f_lw_ARADDR            (arm_a9_hps_h2f_lw_axi_master_araddr),                //                  .araddr
		.h2f_lw_ARLEN             (arm_a9_hps_h2f_lw_axi_master_arlen),                 //                  .arlen
		.h2f_lw_ARSIZE            (arm_a9_hps_h2f_lw_axi_master_arsize),                //                  .arsize
		.h2f_lw_ARBURST           (arm_a9_hps_h2f_lw_axi_master_arburst),               //                  .arburst
		.h2f_lw_ARLOCK            (arm_a9_hps_h2f_lw_axi_master_arlock),                //                  .arlock
		.h2f_lw_ARCACHE           (arm_a9_hps_h2f_lw_axi_master_arcache),               //                  .arcache
		.h2f_lw_ARPROT            (arm_a9_hps_h2f_lw_axi_master_arprot),                //                  .arprot
		.h2f_lw_ARVALID           (arm_a9_hps_h2f_lw_axi_master_arvalid),               //                  .arvalid
		.h2f_lw_ARREADY           (arm_a9_hps_h2f_lw_axi_master_arready),               //                  .arready
		.h2f_lw_RID               (arm_a9_hps_h2f_lw_axi_master_rid),                   //                  .rid
		.h2f_lw_RDATA             (arm_a9_hps_h2f_lw_axi_master_rdata),                 //                  .rdata
		.h2f_lw_RRESP             (arm_a9_hps_h2f_lw_axi_master_rresp),                 //                  .rresp
		.h2f_lw_RLAST             (arm_a9_hps_h2f_lw_axi_master_rlast),                 //                  .rlast
		.h2f_lw_RVALID            (arm_a9_hps_h2f_lw_axi_master_rvalid),                //                  .rvalid
		.h2f_lw_RREADY            (arm_a9_hps_h2f_lw_axi_master_rready),                //                  .rready
		.f2h_irq_p0               (arm_a9_hps_f2h_irq0_irq),                            //          f2h_irq0.irq
		.f2h_irq_p1               (arm_a9_hps_f2h_irq1_irq)                             //          f2h_irq1.irq
	);

	CPEN391_Computer_HEX0_1 hex0_1 (
		.clk        (system_pll_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_hex0_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex0_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex0_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_1_s1_readdata),   //                    .readdata
		.out_port   (hex0_1_export)                           // external_connection.export
	);

	CPEN391_Computer_HEX0_1 hex2_3 (
		.clk        (system_pll_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_hex2_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex2_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex2_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex2_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex2_3_s1_readdata),   //                    .readdata
		.out_port   (hex2_3_export)                           // external_connection.export
	);

	CPEN391_Computer_HEX0_1 hex4_5 (
		.clk        (system_pll_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_hex4_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex4_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex4_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex4_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex4_5_s1_readdata),   //                    .readdata
		.out_port   (hex4_5_export)                           // external_connection.export
	);

	CPEN391_Computer_IO_Bridge io_bridge (
		.clk                (system_pll_sys_clk_clk),                               //                clk.clk
		.reset              (rst_controller_reset_out_reset),                       //              reset.reset
		.avalon_address     (mm_interconnect_0_io_bridge_avalon_slave_address),     //       avalon_slave.address
		.avalon_byteenable  (mm_interconnect_0_io_bridge_avalon_slave_byteenable),  //                   .byteenable
		.avalon_chipselect  (mm_interconnect_0_io_bridge_avalon_slave_chipselect),  //                   .chipselect
		.avalon_read        (mm_interconnect_0_io_bridge_avalon_slave_read),        //                   .read
		.avalon_write       (mm_interconnect_0_io_bridge_avalon_slave_write),       //                   .write
		.avalon_writedata   (mm_interconnect_0_io_bridge_avalon_slave_writedata),   //                   .writedata
		.avalon_readdata    (mm_interconnect_0_io_bridge_avalon_slave_readdata),    //                   .readdata
		.avalon_waitrequest (mm_interconnect_0_io_bridge_avalon_slave_waitrequest), //                   .waitrequest
		.avalon_irq         (irq_mapper_receiver0_irq),                             //          interrupt.irq
		.acknowledge        (io_acknowledge),                                       // external_interface.export
		.irq                (io_irq),                                               //                   .export
		.address            (io_address),                                           //                   .export
		.bus_enable         (io_bus_enable),                                        //                   .export
		.byte_enable        (io_byte_enable),                                       //                   .export
		.rw                 (io_rw),                                                //                   .export
		.write_data         (io_write_data),                                        //                   .export
		.read_data          (io_read_data)                                          //                   .export
	);

	CPEN391_Computer_Interval_Timer interval_timer (
		.clk        (system_pll_sys_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                        //   irq.irq
	);

	CPEN391_Computer_JTAG_To_FPGA_Bridge #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_to_fpga_bridge (
		.clk_clk              (system_pll_sys_clk_clk),                   //          clk.clk
		.clk_reset_reset      (rst_controller_001_reset_out_reset),       //    clk_reset.reset
		.master_address       (jtag_to_fpga_bridge_master_address),       //       master.address
		.master_readdata      (jtag_to_fpga_bridge_master_readdata),      //             .readdata
		.master_read          (jtag_to_fpga_bridge_master_read),          //             .read
		.master_write         (jtag_to_fpga_bridge_master_write),         //             .write
		.master_writedata     (jtag_to_fpga_bridge_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_to_fpga_bridge_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_to_fpga_bridge_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_to_fpga_bridge_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                          // master_reset.reset
	);

	CPEN391_Computer_JTAG_To_FPGA_Bridge #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_to_hps_bridge (
		.clk_clk              (system_pll_sys_clk_clk),                  //          clk.clk
		.clk_reset_reset      (rst_controller_002_reset_out_reset),      //    clk_reset.reset
		.master_address       (jtag_to_hps_bridge_master_address),       //       master.address
		.master_readdata      (jtag_to_hps_bridge_master_readdata),      //             .readdata
		.master_read          (jtag_to_hps_bridge_master_read),          //             .read
		.master_write         (jtag_to_hps_bridge_master_write),         //             .write
		.master_writedata     (jtag_to_hps_bridge_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_to_hps_bridge_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_to_hps_bridge_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_to_hps_bridge_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                         // master_reset.reset
	);

	CPEN391_Computer_JTAG_UART_For_ARM0 jtag_uart_for_arm0 (
		.clk            (system_pll_sys_clk_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                            //               irq.irq
	);

	CPEN391_Computer_JTAG_UART_For_ARM0 jtag_uart_for_arm1 (
		.clk            (system_pll_sys_clk_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver0_irq)                                        //               irq.irq
	);

	CPEN391_Computer_LEDS leds (
		.clk        (system_pll_sys_clk_clk),               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	CPEN391_Computer_Onchip_SRAM onchip_sram (
		.address     (mm_interconnect_0_onchip_sram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_sram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_sram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_sram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_sram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_sram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_sram_s1_byteenable), //       .byteenable
		.address2    (),                                            //     s2.address
		.chipselect2 (),                                            //       .chipselect
		.clken2      (),                                            //       .clken
		.write2      (),                                            //       .write
		.readdata2   (),                                            //       .readdata
		.writedata2  (),                                            //       .writedata
		.byteenable2 (),                                            //       .byteenable
		.clk         (system_pll_sys_clk_clk),                      //   clk1.clk
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	CPEN391_Computer_PushButtons pushbuttons (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pushbuttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pushbuttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pushbuttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pushbuttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pushbuttons_s1_readdata),   //                    .readdata
		.in_port    (pushbuttons_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                     //                 irq.irq
	);

	CPEN391_Computer_SDRAM sdram (
		.clk            (system_pll_sys_clk_clk),                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	CPEN391_Computer_Slider_Switches slider_switches (
		.clk      (system_pll_sys_clk_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_slider_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_slider_switches_s1_readdata), //                    .readdata
		.in_port  (slider_switches_export)                         // external_connection.export
	);

	CPEN391_Computer_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                 //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	render renderer_0 (
		.clk               (system_pll_sys_clk_clk),                         //   clock.clk
		.slave_waitrequest (mm_interconnect_0_renderer_0_slave_waitrequest), //   slave.waitrequest
		.slave_address     (mm_interconnect_0_renderer_0_slave_address),     //        .address
		.slave_read        (mm_interconnect_0_renderer_0_slave_read),        //        .read
		.slave_readdata    (mm_interconnect_0_renderer_0_slave_readdata),    //        .readdata
		.slave_write       (mm_interconnect_0_renderer_0_slave_write),       //        .write
		.slave_writedata   (mm_interconnect_0_renderer_0_slave_writedata),   //        .writedata
		.VGA_R             (vga_vga_r),                                      // conduit.vga_r
		.VGA_G             (vga_vga_g),                                      //        .vga_g
		.VGA_B             (vga_vga_b),                                      //        .vga_b
		.VGA_BLANK_N       (vga_vga_blank_n),                                //        .vga_blank_n
		.VGA_CLK           (vga_vga_clk),                                    //        .vga_clk
		.VGA_HS            (vga_vga_hs),                                     //        .vga_hs
		.VGA_SYNC_N        (vga_vga_sync_n),                                 //        .vga_sync_n
		.VGA_VS            (vga_vga_vs),                                     //        .vga_vs
		.rst_n             (~rst_controller_reset_out_reset)                 //   reset.reset_n
	);

	CPEN391_Computer_sysid_qsys_0 sysid_qsys_0 (
		.clock    (system_pll_sys_clk_clk),                                //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	CPEN391_Computer_mm_interconnect_0 mm_interconnect_0 (
		.ARM_A9_HPS_h2f_axi_master_awid                                        (arm_a9_hps_h2f_axi_master_awid),                                     //                                       ARM_A9_HPS_h2f_axi_master.awid
		.ARM_A9_HPS_h2f_axi_master_awaddr                                      (arm_a9_hps_h2f_axi_master_awaddr),                                   //                                                                .awaddr
		.ARM_A9_HPS_h2f_axi_master_awlen                                       (arm_a9_hps_h2f_axi_master_awlen),                                    //                                                                .awlen
		.ARM_A9_HPS_h2f_axi_master_awsize                                      (arm_a9_hps_h2f_axi_master_awsize),                                   //                                                                .awsize
		.ARM_A9_HPS_h2f_axi_master_awburst                                     (arm_a9_hps_h2f_axi_master_awburst),                                  //                                                                .awburst
		.ARM_A9_HPS_h2f_axi_master_awlock                                      (arm_a9_hps_h2f_axi_master_awlock),                                   //                                                                .awlock
		.ARM_A9_HPS_h2f_axi_master_awcache                                     (arm_a9_hps_h2f_axi_master_awcache),                                  //                                                                .awcache
		.ARM_A9_HPS_h2f_axi_master_awprot                                      (arm_a9_hps_h2f_axi_master_awprot),                                   //                                                                .awprot
		.ARM_A9_HPS_h2f_axi_master_awvalid                                     (arm_a9_hps_h2f_axi_master_awvalid),                                  //                                                                .awvalid
		.ARM_A9_HPS_h2f_axi_master_awready                                     (arm_a9_hps_h2f_axi_master_awready),                                  //                                                                .awready
		.ARM_A9_HPS_h2f_axi_master_wid                                         (arm_a9_hps_h2f_axi_master_wid),                                      //                                                                .wid
		.ARM_A9_HPS_h2f_axi_master_wdata                                       (arm_a9_hps_h2f_axi_master_wdata),                                    //                                                                .wdata
		.ARM_A9_HPS_h2f_axi_master_wstrb                                       (arm_a9_hps_h2f_axi_master_wstrb),                                    //                                                                .wstrb
		.ARM_A9_HPS_h2f_axi_master_wlast                                       (arm_a9_hps_h2f_axi_master_wlast),                                    //                                                                .wlast
		.ARM_A9_HPS_h2f_axi_master_wvalid                                      (arm_a9_hps_h2f_axi_master_wvalid),                                   //                                                                .wvalid
		.ARM_A9_HPS_h2f_axi_master_wready                                      (arm_a9_hps_h2f_axi_master_wready),                                   //                                                                .wready
		.ARM_A9_HPS_h2f_axi_master_bid                                         (arm_a9_hps_h2f_axi_master_bid),                                      //                                                                .bid
		.ARM_A9_HPS_h2f_axi_master_bresp                                       (arm_a9_hps_h2f_axi_master_bresp),                                    //                                                                .bresp
		.ARM_A9_HPS_h2f_axi_master_bvalid                                      (arm_a9_hps_h2f_axi_master_bvalid),                                   //                                                                .bvalid
		.ARM_A9_HPS_h2f_axi_master_bready                                      (arm_a9_hps_h2f_axi_master_bready),                                   //                                                                .bready
		.ARM_A9_HPS_h2f_axi_master_arid                                        (arm_a9_hps_h2f_axi_master_arid),                                     //                                                                .arid
		.ARM_A9_HPS_h2f_axi_master_araddr                                      (arm_a9_hps_h2f_axi_master_araddr),                                   //                                                                .araddr
		.ARM_A9_HPS_h2f_axi_master_arlen                                       (arm_a9_hps_h2f_axi_master_arlen),                                    //                                                                .arlen
		.ARM_A9_HPS_h2f_axi_master_arsize                                      (arm_a9_hps_h2f_axi_master_arsize),                                   //                                                                .arsize
		.ARM_A9_HPS_h2f_axi_master_arburst                                     (arm_a9_hps_h2f_axi_master_arburst),                                  //                                                                .arburst
		.ARM_A9_HPS_h2f_axi_master_arlock                                      (arm_a9_hps_h2f_axi_master_arlock),                                   //                                                                .arlock
		.ARM_A9_HPS_h2f_axi_master_arcache                                     (arm_a9_hps_h2f_axi_master_arcache),                                  //                                                                .arcache
		.ARM_A9_HPS_h2f_axi_master_arprot                                      (arm_a9_hps_h2f_axi_master_arprot),                                   //                                                                .arprot
		.ARM_A9_HPS_h2f_axi_master_arvalid                                     (arm_a9_hps_h2f_axi_master_arvalid),                                  //                                                                .arvalid
		.ARM_A9_HPS_h2f_axi_master_arready                                     (arm_a9_hps_h2f_axi_master_arready),                                  //                                                                .arready
		.ARM_A9_HPS_h2f_axi_master_rid                                         (arm_a9_hps_h2f_axi_master_rid),                                      //                                                                .rid
		.ARM_A9_HPS_h2f_axi_master_rdata                                       (arm_a9_hps_h2f_axi_master_rdata),                                    //                                                                .rdata
		.ARM_A9_HPS_h2f_axi_master_rresp                                       (arm_a9_hps_h2f_axi_master_rresp),                                    //                                                                .rresp
		.ARM_A9_HPS_h2f_axi_master_rlast                                       (arm_a9_hps_h2f_axi_master_rlast),                                    //                                                                .rlast
		.ARM_A9_HPS_h2f_axi_master_rvalid                                      (arm_a9_hps_h2f_axi_master_rvalid),                                   //                                                                .rvalid
		.ARM_A9_HPS_h2f_axi_master_rready                                      (arm_a9_hps_h2f_axi_master_rready),                                   //                                                                .rready
		.ARM_A9_HPS_h2f_lw_axi_master_awid                                     (arm_a9_hps_h2f_lw_axi_master_awid),                                  //                                    ARM_A9_HPS_h2f_lw_axi_master.awid
		.ARM_A9_HPS_h2f_lw_axi_master_awaddr                                   (arm_a9_hps_h2f_lw_axi_master_awaddr),                                //                                                                .awaddr
		.ARM_A9_HPS_h2f_lw_axi_master_awlen                                    (arm_a9_hps_h2f_lw_axi_master_awlen),                                 //                                                                .awlen
		.ARM_A9_HPS_h2f_lw_axi_master_awsize                                   (arm_a9_hps_h2f_lw_axi_master_awsize),                                //                                                                .awsize
		.ARM_A9_HPS_h2f_lw_axi_master_awburst                                  (arm_a9_hps_h2f_lw_axi_master_awburst),                               //                                                                .awburst
		.ARM_A9_HPS_h2f_lw_axi_master_awlock                                   (arm_a9_hps_h2f_lw_axi_master_awlock),                                //                                                                .awlock
		.ARM_A9_HPS_h2f_lw_axi_master_awcache                                  (arm_a9_hps_h2f_lw_axi_master_awcache),                               //                                                                .awcache
		.ARM_A9_HPS_h2f_lw_axi_master_awprot                                   (arm_a9_hps_h2f_lw_axi_master_awprot),                                //                                                                .awprot
		.ARM_A9_HPS_h2f_lw_axi_master_awvalid                                  (arm_a9_hps_h2f_lw_axi_master_awvalid),                               //                                                                .awvalid
		.ARM_A9_HPS_h2f_lw_axi_master_awready                                  (arm_a9_hps_h2f_lw_axi_master_awready),                               //                                                                .awready
		.ARM_A9_HPS_h2f_lw_axi_master_wid                                      (arm_a9_hps_h2f_lw_axi_master_wid),                                   //                                                                .wid
		.ARM_A9_HPS_h2f_lw_axi_master_wdata                                    (arm_a9_hps_h2f_lw_axi_master_wdata),                                 //                                                                .wdata
		.ARM_A9_HPS_h2f_lw_axi_master_wstrb                                    (arm_a9_hps_h2f_lw_axi_master_wstrb),                                 //                                                                .wstrb
		.ARM_A9_HPS_h2f_lw_axi_master_wlast                                    (arm_a9_hps_h2f_lw_axi_master_wlast),                                 //                                                                .wlast
		.ARM_A9_HPS_h2f_lw_axi_master_wvalid                                   (arm_a9_hps_h2f_lw_axi_master_wvalid),                                //                                                                .wvalid
		.ARM_A9_HPS_h2f_lw_axi_master_wready                                   (arm_a9_hps_h2f_lw_axi_master_wready),                                //                                                                .wready
		.ARM_A9_HPS_h2f_lw_axi_master_bid                                      (arm_a9_hps_h2f_lw_axi_master_bid),                                   //                                                                .bid
		.ARM_A9_HPS_h2f_lw_axi_master_bresp                                    (arm_a9_hps_h2f_lw_axi_master_bresp),                                 //                                                                .bresp
		.ARM_A9_HPS_h2f_lw_axi_master_bvalid                                   (arm_a9_hps_h2f_lw_axi_master_bvalid),                                //                                                                .bvalid
		.ARM_A9_HPS_h2f_lw_axi_master_bready                                   (arm_a9_hps_h2f_lw_axi_master_bready),                                //                                                                .bready
		.ARM_A9_HPS_h2f_lw_axi_master_arid                                     (arm_a9_hps_h2f_lw_axi_master_arid),                                  //                                                                .arid
		.ARM_A9_HPS_h2f_lw_axi_master_araddr                                   (arm_a9_hps_h2f_lw_axi_master_araddr),                                //                                                                .araddr
		.ARM_A9_HPS_h2f_lw_axi_master_arlen                                    (arm_a9_hps_h2f_lw_axi_master_arlen),                                 //                                                                .arlen
		.ARM_A9_HPS_h2f_lw_axi_master_arsize                                   (arm_a9_hps_h2f_lw_axi_master_arsize),                                //                                                                .arsize
		.ARM_A9_HPS_h2f_lw_axi_master_arburst                                  (arm_a9_hps_h2f_lw_axi_master_arburst),                               //                                                                .arburst
		.ARM_A9_HPS_h2f_lw_axi_master_arlock                                   (arm_a9_hps_h2f_lw_axi_master_arlock),                                //                                                                .arlock
		.ARM_A9_HPS_h2f_lw_axi_master_arcache                                  (arm_a9_hps_h2f_lw_axi_master_arcache),                               //                                                                .arcache
		.ARM_A9_HPS_h2f_lw_axi_master_arprot                                   (arm_a9_hps_h2f_lw_axi_master_arprot),                                //                                                                .arprot
		.ARM_A9_HPS_h2f_lw_axi_master_arvalid                                  (arm_a9_hps_h2f_lw_axi_master_arvalid),                               //                                                                .arvalid
		.ARM_A9_HPS_h2f_lw_axi_master_arready                                  (arm_a9_hps_h2f_lw_axi_master_arready),                               //                                                                .arready
		.ARM_A9_HPS_h2f_lw_axi_master_rid                                      (arm_a9_hps_h2f_lw_axi_master_rid),                                   //                                                                .rid
		.ARM_A9_HPS_h2f_lw_axi_master_rdata                                    (arm_a9_hps_h2f_lw_axi_master_rdata),                                 //                                                                .rdata
		.ARM_A9_HPS_h2f_lw_axi_master_rresp                                    (arm_a9_hps_h2f_lw_axi_master_rresp),                                 //                                                                .rresp
		.ARM_A9_HPS_h2f_lw_axi_master_rlast                                    (arm_a9_hps_h2f_lw_axi_master_rlast),                                 //                                                                .rlast
		.ARM_A9_HPS_h2f_lw_axi_master_rvalid                                   (arm_a9_hps_h2f_lw_axi_master_rvalid),                                //                                                                .rvalid
		.ARM_A9_HPS_h2f_lw_axi_master_rready                                   (arm_a9_hps_h2f_lw_axi_master_rready),                                //                                                                .rready
		.System_PLL_sys_clk_clk                                                (system_pll_sys_clk_clk),                                             //                                              System_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                                 // ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.JTAG_To_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                     //             JTAG_To_FPGA_Bridge_clk_reset_reset_bridge_in_reset.reset
		.SDRAM_reset_reset_bridge_in_reset_reset                               (rst_controller_reset_out_reset),                                     //                               SDRAM_reset_reset_bridge_in_reset.reset
		.JTAG_To_FPGA_Bridge_master_address                                    (jtag_to_fpga_bridge_master_address),                                 //                                      JTAG_To_FPGA_Bridge_master.address
		.JTAG_To_FPGA_Bridge_master_waitrequest                                (jtag_to_fpga_bridge_master_waitrequest),                             //                                                                .waitrequest
		.JTAG_To_FPGA_Bridge_master_byteenable                                 (jtag_to_fpga_bridge_master_byteenable),                              //                                                                .byteenable
		.JTAG_To_FPGA_Bridge_master_read                                       (jtag_to_fpga_bridge_master_read),                                    //                                                                .read
		.JTAG_To_FPGA_Bridge_master_readdata                                   (jtag_to_fpga_bridge_master_readdata),                                //                                                                .readdata
		.JTAG_To_FPGA_Bridge_master_readdatavalid                              (jtag_to_fpga_bridge_master_readdatavalid),                           //                                                                .readdatavalid
		.JTAG_To_FPGA_Bridge_master_write                                      (jtag_to_fpga_bridge_master_write),                                   //                                                                .write
		.JTAG_To_FPGA_Bridge_master_writedata                                  (jtag_to_fpga_bridge_master_writedata),                               //                                                                .writedata
		.HEX0_1_s1_address                                                     (mm_interconnect_0_hex0_1_s1_address),                                //                                                       HEX0_1_s1.address
		.HEX0_1_s1_write                                                       (mm_interconnect_0_hex0_1_s1_write),                                  //                                                                .write
		.HEX0_1_s1_readdata                                                    (mm_interconnect_0_hex0_1_s1_readdata),                               //                                                                .readdata
		.HEX0_1_s1_writedata                                                   (mm_interconnect_0_hex0_1_s1_writedata),                              //                                                                .writedata
		.HEX0_1_s1_chipselect                                                  (mm_interconnect_0_hex0_1_s1_chipselect),                             //                                                                .chipselect
		.HEX2_3_s1_address                                                     (mm_interconnect_0_hex2_3_s1_address),                                //                                                       HEX2_3_s1.address
		.HEX2_3_s1_write                                                       (mm_interconnect_0_hex2_3_s1_write),                                  //                                                                .write
		.HEX2_3_s1_readdata                                                    (mm_interconnect_0_hex2_3_s1_readdata),                               //                                                                .readdata
		.HEX2_3_s1_writedata                                                   (mm_interconnect_0_hex2_3_s1_writedata),                              //                                                                .writedata
		.HEX2_3_s1_chipselect                                                  (mm_interconnect_0_hex2_3_s1_chipselect),                             //                                                                .chipselect
		.HEX4_5_s1_address                                                     (mm_interconnect_0_hex4_5_s1_address),                                //                                                       HEX4_5_s1.address
		.HEX4_5_s1_write                                                       (mm_interconnect_0_hex4_5_s1_write),                                  //                                                                .write
		.HEX4_5_s1_readdata                                                    (mm_interconnect_0_hex4_5_s1_readdata),                               //                                                                .readdata
		.HEX4_5_s1_writedata                                                   (mm_interconnect_0_hex4_5_s1_writedata),                              //                                                                .writedata
		.HEX4_5_s1_chipselect                                                  (mm_interconnect_0_hex4_5_s1_chipselect),                             //                                                                .chipselect
		.Interval_Timer_s1_address                                             (mm_interconnect_0_interval_timer_s1_address),                        //                                               Interval_Timer_s1.address
		.Interval_Timer_s1_write                                               (mm_interconnect_0_interval_timer_s1_write),                          //                                                                .write
		.Interval_Timer_s1_readdata                                            (mm_interconnect_0_interval_timer_s1_readdata),                       //                                                                .readdata
		.Interval_Timer_s1_writedata                                           (mm_interconnect_0_interval_timer_s1_writedata),                      //                                                                .writedata
		.Interval_Timer_s1_chipselect                                          (mm_interconnect_0_interval_timer_s1_chipselect),                     //                                                                .chipselect
		.IO_Bridge_avalon_slave_address                                        (mm_interconnect_0_io_bridge_avalon_slave_address),                   //                                          IO_Bridge_avalon_slave.address
		.IO_Bridge_avalon_slave_write                                          (mm_interconnect_0_io_bridge_avalon_slave_write),                     //                                                                .write
		.IO_Bridge_avalon_slave_read                                           (mm_interconnect_0_io_bridge_avalon_slave_read),                      //                                                                .read
		.IO_Bridge_avalon_slave_readdata                                       (mm_interconnect_0_io_bridge_avalon_slave_readdata),                  //                                                                .readdata
		.IO_Bridge_avalon_slave_writedata                                      (mm_interconnect_0_io_bridge_avalon_slave_writedata),                 //                                                                .writedata
		.IO_Bridge_avalon_slave_byteenable                                     (mm_interconnect_0_io_bridge_avalon_slave_byteenable),                //                                                                .byteenable
		.IO_Bridge_avalon_slave_waitrequest                                    (mm_interconnect_0_io_bridge_avalon_slave_waitrequest),               //                                                                .waitrequest
		.IO_Bridge_avalon_slave_chipselect                                     (mm_interconnect_0_io_bridge_avalon_slave_chipselect),                //                                                                .chipselect
		.JTAG_UART_For_ARM0_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_address),     //                            JTAG_UART_For_ARM0_avalon_jtag_slave.address
		.JTAG_UART_For_ARM0_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_write),       //                                                                .write
		.JTAG_UART_For_ARM0_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_read),        //                                                                .read
		.JTAG_UART_For_ARM0_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_readdata),    //                                                                .readdata
		.JTAG_UART_For_ARM0_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_writedata),   //                                                                .writedata
		.JTAG_UART_For_ARM0_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_waitrequest), //                                                                .waitrequest
		.JTAG_UART_For_ARM0_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_for_arm0_avalon_jtag_slave_chipselect),  //                                                                .chipselect
		.JTAG_UART_For_ARM1_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_address),     //                            JTAG_UART_For_ARM1_avalon_jtag_slave.address
		.JTAG_UART_For_ARM1_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_write),       //                                                                .write
		.JTAG_UART_For_ARM1_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_read),        //                                                                .read
		.JTAG_UART_For_ARM1_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_readdata),    //                                                                .readdata
		.JTAG_UART_For_ARM1_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_writedata),   //                                                                .writedata
		.JTAG_UART_For_ARM1_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_waitrequest), //                                                                .waitrequest
		.JTAG_UART_For_ARM1_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_for_arm1_avalon_jtag_slave_chipselect),  //                                                                .chipselect
		.LEDS_s1_address                                                       (mm_interconnect_0_leds_s1_address),                                  //                                                         LEDS_s1.address
		.LEDS_s1_write                                                         (mm_interconnect_0_leds_s1_write),                                    //                                                                .write
		.LEDS_s1_readdata                                                      (mm_interconnect_0_leds_s1_readdata),                                 //                                                                .readdata
		.LEDS_s1_writedata                                                     (mm_interconnect_0_leds_s1_writedata),                                //                                                                .writedata
		.LEDS_s1_chipselect                                                    (mm_interconnect_0_leds_s1_chipselect),                               //                                                                .chipselect
		.Onchip_SRAM_s1_address                                                (mm_interconnect_0_onchip_sram_s1_address),                           //                                                  Onchip_SRAM_s1.address
		.Onchip_SRAM_s1_write                                                  (mm_interconnect_0_onchip_sram_s1_write),                             //                                                                .write
		.Onchip_SRAM_s1_readdata                                               (mm_interconnect_0_onchip_sram_s1_readdata),                          //                                                                .readdata
		.Onchip_SRAM_s1_writedata                                              (mm_interconnect_0_onchip_sram_s1_writedata),                         //                                                                .writedata
		.Onchip_SRAM_s1_byteenable                                             (mm_interconnect_0_onchip_sram_s1_byteenable),                        //                                                                .byteenable
		.Onchip_SRAM_s1_chipselect                                             (mm_interconnect_0_onchip_sram_s1_chipselect),                        //                                                                .chipselect
		.Onchip_SRAM_s1_clken                                                  (mm_interconnect_0_onchip_sram_s1_clken),                             //                                                                .clken
		.PushButtons_s1_address                                                (mm_interconnect_0_pushbuttons_s1_address),                           //                                                  PushButtons_s1.address
		.PushButtons_s1_write                                                  (mm_interconnect_0_pushbuttons_s1_write),                             //                                                                .write
		.PushButtons_s1_readdata                                               (mm_interconnect_0_pushbuttons_s1_readdata),                          //                                                                .readdata
		.PushButtons_s1_writedata                                              (mm_interconnect_0_pushbuttons_s1_writedata),                         //                                                                .writedata
		.PushButtons_s1_chipselect                                             (mm_interconnect_0_pushbuttons_s1_chipselect),                        //                                                                .chipselect
		.renderer_0_slave_address                                              (mm_interconnect_0_renderer_0_slave_address),                         //                                                renderer_0_slave.address
		.renderer_0_slave_write                                                (mm_interconnect_0_renderer_0_slave_write),                           //                                                                .write
		.renderer_0_slave_read                                                 (mm_interconnect_0_renderer_0_slave_read),                            //                                                                .read
		.renderer_0_slave_readdata                                             (mm_interconnect_0_renderer_0_slave_readdata),                        //                                                                .readdata
		.renderer_0_slave_writedata                                            (mm_interconnect_0_renderer_0_slave_writedata),                       //                                                                .writedata
		.renderer_0_slave_waitrequest                                          (mm_interconnect_0_renderer_0_slave_waitrequest),                     //                                                                .waitrequest
		.SDRAM_s1_address                                                      (mm_interconnect_0_sdram_s1_address),                                 //                                                        SDRAM_s1.address
		.SDRAM_s1_write                                                        (mm_interconnect_0_sdram_s1_write),                                   //                                                                .write
		.SDRAM_s1_read                                                         (mm_interconnect_0_sdram_s1_read),                                    //                                                                .read
		.SDRAM_s1_readdata                                                     (mm_interconnect_0_sdram_s1_readdata),                                //                                                                .readdata
		.SDRAM_s1_writedata                                                    (mm_interconnect_0_sdram_s1_writedata),                               //                                                                .writedata
		.SDRAM_s1_byteenable                                                   (mm_interconnect_0_sdram_s1_byteenable),                              //                                                                .byteenable
		.SDRAM_s1_readdatavalid                                                (mm_interconnect_0_sdram_s1_readdatavalid),                           //                                                                .readdatavalid
		.SDRAM_s1_waitrequest                                                  (mm_interconnect_0_sdram_s1_waitrequest),                             //                                                                .waitrequest
		.SDRAM_s1_chipselect                                                   (mm_interconnect_0_sdram_s1_chipselect),                              //                                                                .chipselect
		.Slider_Switches_s1_address                                            (mm_interconnect_0_slider_switches_s1_address),                       //                                              Slider_Switches_s1.address
		.Slider_Switches_s1_readdata                                           (mm_interconnect_0_slider_switches_s1_readdata),                      //                                                                .readdata
		.sysid_qsys_0_control_slave_address                                    (mm_interconnect_0_sysid_qsys_0_control_slave_address),               //                                      sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                                   (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)               //                                                                .readdata
	);

	CPEN391_Computer_mm_interconnect_1 mm_interconnect_1 (
		.ARM_A9_HPS_f2h_axi_slave_awid                                          (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid),    //                                         ARM_A9_HPS_f2h_axi_slave.awid
		.ARM_A9_HPS_f2h_axi_slave_awaddr                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr),  //                                                                 .awaddr
		.ARM_A9_HPS_f2h_axi_slave_awlen                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen),   //                                                                 .awlen
		.ARM_A9_HPS_f2h_axi_slave_awsize                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize),  //                                                                 .awsize
		.ARM_A9_HPS_f2h_axi_slave_awburst                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst), //                                                                 .awburst
		.ARM_A9_HPS_f2h_axi_slave_awlock                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock),  //                                                                 .awlock
		.ARM_A9_HPS_f2h_axi_slave_awcache                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache), //                                                                 .awcache
		.ARM_A9_HPS_f2h_axi_slave_awprot                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot),  //                                                                 .awprot
		.ARM_A9_HPS_f2h_axi_slave_awuser                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser),  //                                                                 .awuser
		.ARM_A9_HPS_f2h_axi_slave_awvalid                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid), //                                                                 .awvalid
		.ARM_A9_HPS_f2h_axi_slave_awready                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready), //                                                                 .awready
		.ARM_A9_HPS_f2h_axi_slave_wid                                           (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid),     //                                                                 .wid
		.ARM_A9_HPS_f2h_axi_slave_wdata                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata),   //                                                                 .wdata
		.ARM_A9_HPS_f2h_axi_slave_wstrb                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb),   //                                                                 .wstrb
		.ARM_A9_HPS_f2h_axi_slave_wlast                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast),   //                                                                 .wlast
		.ARM_A9_HPS_f2h_axi_slave_wvalid                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid),  //                                                                 .wvalid
		.ARM_A9_HPS_f2h_axi_slave_wready                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready),  //                                                                 .wready
		.ARM_A9_HPS_f2h_axi_slave_bid                                           (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid),     //                                                                 .bid
		.ARM_A9_HPS_f2h_axi_slave_bresp                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp),   //                                                                 .bresp
		.ARM_A9_HPS_f2h_axi_slave_bvalid                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid),  //                                                                 .bvalid
		.ARM_A9_HPS_f2h_axi_slave_bready                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready),  //                                                                 .bready
		.ARM_A9_HPS_f2h_axi_slave_arid                                          (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid),    //                                                                 .arid
		.ARM_A9_HPS_f2h_axi_slave_araddr                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr),  //                                                                 .araddr
		.ARM_A9_HPS_f2h_axi_slave_arlen                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen),   //                                                                 .arlen
		.ARM_A9_HPS_f2h_axi_slave_arsize                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize),  //                                                                 .arsize
		.ARM_A9_HPS_f2h_axi_slave_arburst                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst), //                                                                 .arburst
		.ARM_A9_HPS_f2h_axi_slave_arlock                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock),  //                                                                 .arlock
		.ARM_A9_HPS_f2h_axi_slave_arcache                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache), //                                                                 .arcache
		.ARM_A9_HPS_f2h_axi_slave_arprot                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot),  //                                                                 .arprot
		.ARM_A9_HPS_f2h_axi_slave_aruser                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser),  //                                                                 .aruser
		.ARM_A9_HPS_f2h_axi_slave_arvalid                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid), //                                                                 .arvalid
		.ARM_A9_HPS_f2h_axi_slave_arready                                       (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready), //                                                                 .arready
		.ARM_A9_HPS_f2h_axi_slave_rid                                           (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid),     //                                                                 .rid
		.ARM_A9_HPS_f2h_axi_slave_rdata                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata),   //                                                                 .rdata
		.ARM_A9_HPS_f2h_axi_slave_rresp                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp),   //                                                                 .rresp
		.ARM_A9_HPS_f2h_axi_slave_rlast                                         (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast),   //                                                                 .rlast
		.ARM_A9_HPS_f2h_axi_slave_rvalid                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid),  //                                                                 .rvalid
		.ARM_A9_HPS_f2h_axi_slave_rready                                        (mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready),  //                                                                 .rready
		.System_PLL_sys_clk_clk                                                 (system_pll_sys_clk_clk),                             //                                               System_PLL_sys_clk.clk
		.ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset  (rst_controller_003_reset_out_reset),                 //  ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.JTAG_To_HPS_Bridge_clk_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                     //               JTAG_To_HPS_Bridge_clk_reset_reset_bridge_in_reset.reset
		.JTAG_To_HPS_Bridge_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                     // JTAG_To_HPS_Bridge_master_translator_reset_reset_bridge_in_reset.reset
		.JTAG_To_HPS_Bridge_master_address                                      (jtag_to_hps_bridge_master_address),                  //                                        JTAG_To_HPS_Bridge_master.address
		.JTAG_To_HPS_Bridge_master_waitrequest                                  (jtag_to_hps_bridge_master_waitrequest),              //                                                                 .waitrequest
		.JTAG_To_HPS_Bridge_master_byteenable                                   (jtag_to_hps_bridge_master_byteenable),               //                                                                 .byteenable
		.JTAG_To_HPS_Bridge_master_read                                         (jtag_to_hps_bridge_master_read),                     //                                                                 .read
		.JTAG_To_HPS_Bridge_master_readdata                                     (jtag_to_hps_bridge_master_readdata),                 //                                                                 .readdata
		.JTAG_To_HPS_Bridge_master_readdatavalid                                (jtag_to_hps_bridge_master_readdatavalid),            //                                                                 .readdatavalid
		.JTAG_To_HPS_Bridge_master_write                                        (jtag_to_hps_bridge_master_write),                    //                                                                 .write
		.JTAG_To_HPS_Bridge_master_writedata                                    (jtag_to_hps_bridge_master_writedata)                 //                                                                 .writedata
	);

	CPEN391_Computer_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq), // receiver3.irq
		.sender_irq    (arm_a9_hps_f2h_irq0_irq)   //    sender.irq
	);

	CPEN391_Computer_irq_mapper_001 irq_mapper_001 (
		.clk           (),                             //       clk.clk
		.reset         (),                             // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq), // receiver0.irq
		.sender_irq    (arm_a9_hps_f2h_irq1_irq)       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
